class core_ibex_vseqr extends uvm_sequencer;

  ibex_mem_intf_response_sequencer                   data_if_seqr;
  ibex_mem_intf_response_sequencer                   instr_if_seqr;

  `uvm_component_utils(core_ibex_vseqr)
  `uvm_component_new

endclass
